LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY toggle_flip_flop IS
    PORT(

    );
END toggle_flip_flop;